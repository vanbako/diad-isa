`ifndef SR_VH
`define SR_VH

`define INDEX_FL  4'h0
`define INDEX_LR  4'h1
`define INDEX_IR  4'h2
`define INDEX_SSP 4'h3
`define INDEX_PC  4'hF

`endif